`timescale 1ns / 1ps
module test_rom
	(
		input wire clk,
		input wire [4:0] row,
		input wire [3:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [3:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		9'b000000000: color_data = 12'b111111111111;
		9'b000000001: color_data = 12'b000000000000;
		9'b000000010: color_data = 12'b000000000000;
		9'b000000011: color_data = 12'b000000000000;
		9'b000000100: color_data = 12'b000000000000;
		9'b000000101: color_data = 12'b000000000000;
		9'b000000110: color_data = 12'b000000000000;
		9'b000000111: color_data = 12'b000000000000;
		9'b000001000: color_data = 12'b000000000000;
		9'b000001001: color_data = 12'b000000000000;

		9'b000010000: color_data = 12'b111111111111;
		9'b000010001: color_data = 12'b000000000000;
		9'b000010010: color_data = 12'b111111111111;
		9'b000010011: color_data = 12'b000000000000;
		9'b000010100: color_data = 12'b000000000000;
		9'b000010101: color_data = 12'b000000000000;
		9'b000010110: color_data = 12'b000000000000;
		9'b000010111: color_data = 12'b000000000000;
		9'b000011000: color_data = 12'b000000000000;
		9'b000011001: color_data = 12'b000000000000;

		9'b000100000: color_data = 12'b000000000000;
		9'b000100001: color_data = 12'b000000000000;
		9'b000100010: color_data = 12'b000000000000;
		9'b000100011: color_data = 12'b000000000000;
		9'b000100100: color_data = 12'b000000000000;
		9'b000100101: color_data = 12'b000000000000;
		9'b000100110: color_data = 12'b000000000000;
		9'b000100111: color_data = 12'b000000000000;
		9'b000101000: color_data = 12'b000000000000;
		9'b000101001: color_data = 12'b000000000000;

		9'b000110000: color_data = 12'b000000000000;
		9'b000110001: color_data = 12'b111111111111;
		9'b000110010: color_data = 12'b111111111111;
		9'b000110011: color_data = 12'b111111111111;
		9'b000110100: color_data = 12'b111111111111;
		9'b000110101: color_data = 12'b111111111111;
		9'b000110110: color_data = 12'b111111111111;
		9'b000110111: color_data = 12'b111111111111;
		9'b000111000: color_data = 12'b111111111111;
		9'b000111001: color_data = 12'b000000000000;

		9'b001000000: color_data = 12'b000000000000;
		9'b001000001: color_data = 12'b111111111111;
		9'b001000010: color_data = 12'b111111111111;
		9'b001000011: color_data = 12'b000000000000;
		9'b001000100: color_data = 12'b111111111111;
		9'b001000101: color_data = 12'b111111111111;
		9'b001000110: color_data = 12'b000000000000;
		9'b001000111: color_data = 12'b111111111111;
		9'b001001000: color_data = 12'b111111111111;
		9'b001001001: color_data = 12'b000000000000;

		9'b001010000: color_data = 12'b000000000000;
		9'b001010001: color_data = 12'b111111111111;
		9'b001010010: color_data = 12'b111111111111;
		9'b001010011: color_data = 12'b111111111111;
		9'b001010100: color_data = 12'b111111111111;
		9'b001010101: color_data = 12'b111111111111;
		9'b001010110: color_data = 12'b111111111111;
		9'b001010111: color_data = 12'b111111111111;
		9'b001011000: color_data = 12'b111111111111;
		9'b001011001: color_data = 12'b000000000000;

		9'b001100000: color_data = 12'b000000000000;
		9'b001100001: color_data = 12'b111111111111;
		9'b001100010: color_data = 12'b111111111111;
		9'b001100011: color_data = 12'b111111111111;
		9'b001100100: color_data = 12'b111111111111;
		9'b001100101: color_data = 12'b111111111111;
		9'b001100110: color_data = 12'b111111111111;
		9'b001100111: color_data = 12'b111111111111;
		9'b001101000: color_data = 12'b111111111111;
		9'b001101001: color_data = 12'b000000000000;

		9'b001110000: color_data = 12'b000000000000;
		9'b001110001: color_data = 12'b000000000000;
		9'b001110010: color_data = 12'b111010001000;
		9'b001110011: color_data = 12'b111111111111;
		9'b001110100: color_data = 12'b111111111111;
		9'b001110101: color_data = 12'b111111111111;
		9'b001110110: color_data = 12'b111010001000;
		9'b001110111: color_data = 12'b111111111111;
		9'b001111000: color_data = 12'b000000000000;
		9'b001111001: color_data = 12'b000000000000;

		9'b010000000: color_data = 12'b000000000000;
		9'b010000001: color_data = 12'b000000000000;
		9'b010000010: color_data = 12'b111010001000;
		9'b010000011: color_data = 12'b111111111111;
		9'b010000100: color_data = 12'b111111111111;
		9'b010000101: color_data = 12'b111111111111;
		9'b010000110: color_data = 12'b111010001000;
		9'b010000111: color_data = 12'b111111111111;
		9'b010001000: color_data = 12'b000000000000;
		9'b010001001: color_data = 12'b000000000000;

		9'b010010000: color_data = 12'b000000000000;
		9'b010010001: color_data = 12'b000000000000;
		9'b010010010: color_data = 12'b111111111111;
		9'b010010011: color_data = 12'b111111111111;
		9'b010010100: color_data = 12'b111111111111;
		9'b010010101: color_data = 12'b111111111111;
		9'b010010110: color_data = 12'b111111111111;
		9'b010010111: color_data = 12'b000000000000;
		9'b010011000: color_data = 12'b000000000000;
		9'b010011001: color_data = 12'b000000000000;

		9'b010100000: color_data = 12'b000000000000;
		9'b010100001: color_data = 12'b000000000000;
		9'b010100010: color_data = 12'b111010001000;
		9'b010100011: color_data = 12'b111111111111;
		9'b010100100: color_data = 12'b111111111111;
		9'b010100101: color_data = 12'b111111111111;
		9'b010100110: color_data = 12'b111010001000;
		9'b010100111: color_data = 12'b000000000000;
		9'b010101000: color_data = 12'b000000000000;
		9'b010101001: color_data = 12'b000000000000;

		9'b010110000: color_data = 12'b000000000000;
		9'b010110001: color_data = 12'b000000000000;
		9'b010110010: color_data = 12'b111111111111;
		9'b010110011: color_data = 12'b111111111111;
		9'b010110100: color_data = 12'b111111111111;
		9'b010110101: color_data = 12'b111111111111;
		9'b010110110: color_data = 12'b000000000000;
		9'b010110111: color_data = 12'b000000000000;
		9'b010111000: color_data = 12'b000000000000;
		9'b010111001: color_data = 12'b000000000000;

		9'b011000000: color_data = 12'b000000000000;
		9'b011000001: color_data = 12'b000000000000;
		9'b011000010: color_data = 12'b000000000000;
		9'b011000011: color_data = 12'b111111111111;
		9'b011000100: color_data = 12'b000000000000;
		9'b011000101: color_data = 12'b111111111111;
		9'b011000110: color_data = 12'b000000000000;
		9'b011000111: color_data = 12'b000000000000;
		9'b011001000: color_data = 12'b000000000000;
		9'b011001001: color_data = 12'b000000000000;

		9'b011010000: color_data = 12'b000000000000;
		9'b011010001: color_data = 12'b000000000000;
		9'b011010010: color_data = 12'b111111111111;
		9'b011010011: color_data = 12'b111111111111;
		9'b011010100: color_data = 12'b111111111111;
		9'b011010101: color_data = 12'b111111111111;
		9'b011010110: color_data = 12'b000000000000;
		9'b011010111: color_data = 12'b000000000000;
		9'b011011000: color_data = 12'b000000000000;
		9'b011011001: color_data = 12'b000000000000;

		9'b011100000: color_data = 12'b000000000000;
		9'b011100001: color_data = 12'b000000000000;
		9'b011100010: color_data = 12'b111111111111;
		9'b011100011: color_data = 12'b111111111111;
		9'b011100100: color_data = 12'b111111111111;
		9'b011100101: color_data = 12'b000000000000;
		9'b011100110: color_data = 12'b000000000000;
		9'b011100111: color_data = 12'b000000000000;
		9'b011101000: color_data = 12'b000000000000;
		9'b011101001: color_data = 12'b000000000000;

		9'b011110000: color_data = 12'b000000000000;
		9'b011110001: color_data = 12'b000000000000;
		9'b011110010: color_data = 12'b000000000000;
		9'b011110011: color_data = 12'b111111111111;
		9'b011110100: color_data = 12'b111111111111;
		9'b011110101: color_data = 12'b000000000000;
		9'b011110110: color_data = 12'b000000000000;
		9'b011110111: color_data = 12'b000000000000;
		9'b011111000: color_data = 12'b000000000000;
		9'b011111001: color_data = 12'b000000000000;

		9'b100000000: color_data = 12'b000000000000;
		9'b100000001: color_data = 12'b000000000000;
		9'b100000010: color_data = 12'b000000000000;
		9'b100000011: color_data = 12'b111111111111;
		9'b100000100: color_data = 12'b000000000000;
		9'b100000101: color_data = 12'b000000000000;
		9'b100000110: color_data = 12'b000000000000;
		9'b100000111: color_data = 12'b000000000000;
		9'b100001000: color_data = 12'b000000000000;
		9'b100001001: color_data = 12'b000000000000;

		9'b100010000: color_data = 12'b000000000000;
		9'b100010001: color_data = 12'b000000000000;
		9'b100010010: color_data = 12'b000000000000;
		9'b100010011: color_data = 12'b111111111111;
		9'b100010100: color_data = 12'b000000000000;
		9'b100010101: color_data = 12'b000000000000;
		9'b100010110: color_data = 12'b000000000000;
		9'b100010111: color_data = 12'b000000000000;
		9'b100011000: color_data = 12'b000000000000;
		9'b100011001: color_data = 12'b000000000000;

		9'b100100000: color_data = 12'b000000000000;
		9'b100100001: color_data = 12'b000000000000;
		9'b100100010: color_data = 12'b000000000000;
		9'b100100011: color_data = 12'b111111111111;
		9'b100100100: color_data = 12'b000000000000;
		9'b100100101: color_data = 12'b000000000000;
		9'b100100110: color_data = 12'b000000000000;
		9'b100100111: color_data = 12'b000000000000;
		9'b100101000: color_data = 12'b000000000000;
		9'b100101001: color_data = 12'b000000000000;

		9'b100110000: color_data = 12'b000000000000;
		9'b100110001: color_data = 12'b000000000000;
		9'b100110010: color_data = 12'b000000000000;
		9'b100110011: color_data = 12'b000000000000;
		9'b100110100: color_data = 12'b000000000000;
		9'b100110101: color_data = 12'b000000000000;
		9'b100110110: color_data = 12'b000000000000;
		9'b100110111: color_data = 12'b000000000000;
		9'b100111000: color_data = 12'b000000000000;
		9'b100111001: color_data = 12'b000000000000;

		default: color_data = 12'b000000000000;
	endcase
endmodule
